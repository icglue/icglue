<%
    ##  icglue - module template
-%>
<%I header.module.template.v %>
<%
    ###########################################
    ## <regfile>
-%>
<%I regfile.module.template.v %>
<%
    ## </regfile>
    ###########################################
-%>

endmodule

<%- # vim: set filetype=verilog_template: -%>
